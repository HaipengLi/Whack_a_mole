

 
 
 

 



window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /hit_mouse_tb/status
      waveform add -signals /hit_mouse_tb/hit_mouse_synth_inst/bmg_port/CLKA
      waveform add -signals /hit_mouse_tb/hit_mouse_synth_inst/bmg_port/ADDRA
      waveform add -signals /hit_mouse_tb/hit_mouse_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
